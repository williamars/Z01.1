corsi@corsi-note.18581:1585446834